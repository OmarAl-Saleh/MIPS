module INST_MEM #(
  parameter size = 10000,          
  parameter data_width = 32    
)(
 // input clk,
  input reset,                   
  input [31:0] address,
  output reg [31:0] inst_out

);
   reg [31:0] inst_mem [0:size - 1];

  
 
integer i ; 

//  endmodule 

reg state = 1'b0;
  
  
//  
  always @(*) 

 begin
        case (state)
            1'b0: begin
                state <= 1'b1;
					 // Enter here the Instructions of the program
					 
					 for (i = 0; i < 2600; i = i + 26) begin
		  //Benchmark 2
		  
			inst_mem[0+i]=32'b00001100000000000000000000000010;
			
			//inst_mem[1+i]=32'b00001000000000000000000000011001; // JUMP End 
			
			inst_mem[1+i]=32'b00010000000000000000000000010111; // beq r0,r0,End (23 instruction between (offset))
			
			inst_mem[2+i]=32'b00100000000100000000000000000000;
			inst_mem[3+i]=32'b00100000000010000000000000000000;
			inst_mem[4+i]=32'b00100000000100010000000000010011;
			inst_mem[5+i]=32'b00011001000100010000000000010010;//sel1
			inst_mem[6+i]=32'b00100000000010010000000000000000;
			inst_mem[7+i]=32'b00000010001010010101000000100010;
			inst_mem[8+i]=32'b00011001001010100000000000001101; // sel2
			inst_mem[9+i]=32'b00000001001000000101100010000000;
			inst_mem[10+i]=32'b00000010000010110110000000100000;
			inst_mem[11+i]=32'b10001101100011010000000000000000;
			inst_mem[12+i]=32'b10001101100011100000000000000100;
			inst_mem[13+i]=32'b00011001101011100000000000000001;
			
		//	inst_mem[14+i]=32'b00001000000000000000000000010100; // Jump --> ES
		
			inst_mem[14+i]=32'b00010000000000000000000000000101;//beq r0,r0,ES (offset 5)
			
			inst_mem[15+i]=32'b00000001101000000111100000100000;
			inst_mem[16+i]=32'b00000001110000000110100000100000;
			inst_mem[17+i]=32'b00000001111000000111000000100000;
			inst_mem[18+i]=32'b10101101100011010000000000000000;
			inst_mem[19+i]=32'b10101101100011100000000000000100;
			inst_mem[20+i]=32'b00100001001010010000000000000001; //ES
			
			//inst_mem[21+i]=32'b00001000000000000000000000001000;//Jump -->  8 sel2
			 
			 inst_mem[21+i]=32'b00010000000000001111111111110010; // beq r0,r0 , sel2 offset(-14)

			
			inst_mem[22+i]=32'b00100001000010000000000000000001;
			
			
		//	inst_mem[23+i]=32'b00001000000000000000000000000101;// JUMP --> 5 sel 1
		
		   inst_mem[23+i]=32'b 00010000000000001111111111101101; // beq r0,r0,sel1 offset(-19)
			
			inst_mem[24+i]=32'b00000011111001010010000000001000;
			inst_mem[25+i]=32'b00000000000000000000000000100000;
	
		
      end
		
	//	beq r0, r0, P1			000100 00000 00000 0000000000000001
					 
//B.2
//inst_mem[0]=32'b00001100000000000000000000000010;
//inst_mem[1]=32'b00001000000000000000000000011001;
//inst_mem[2]=32'b00100000000100000000000000000000;
//inst_mem[3]=32'b00100000000010000000000000000000;
//inst_mem[4]=32'b00100000000100010000000000010011;
//inst_mem[5]=32'b00011001000100010000000000010010;
//inst_mem[6]=32'b00100000000010010000000000000000;
//inst_mem[7]=32'b00000010001010010101000000100010;
//inst_mem[8]=32'b00011001001010100000000000001101;
//inst_mem[9]=32'b00000001001000000101100010000000;
//inst_mem[10]=32'b00000010000010110110000000100000;
//inst_mem[11]=32'b10001101100011010000000000000000;
//inst_mem[12]=32'b10001101100011100000000000000100;
//inst_mem[13]=32'b00011001101011100000000000000001;
//inst_mem[14]=32'b00001000000000000000000000010100;
//inst_mem[15]=32'b00000001101000000111100000100000;
//inst_mem[16]=32'b00000001110000000110100000100000;
//inst_mem[17]=32'b00000001111000000111000000100000;
//inst_mem[18]=32'b10101101100011010000000000000000;
//inst_mem[19]=32'b10101101100011100000000000000100;
//inst_mem[20]=32'b00100001001010010000000000000001;
//inst_mem[21]=32'b00001000000000000000000000001000;
//inst_mem[22]=32'b00100001000010000000000000000001;
//inst_mem[23]=32'b00001000000000000000000000000101;
//inst_mem[24]=32'b00000011111001010010000000001000;
//inst_mem[25]=32'b00000000000000000000000000100000;
					 
					 //B.1

//inst_mem[0]=32'b10001100000000010000000000000000;
//inst_mem[1]=32'b00110100000000100000000000000100;
//inst_mem[2]=32'b00100000000000111111111111111110;
//inst_mem[3]=32'b10001100000001000000000000000100;
//inst_mem[4]=32'b00000000001000010010100000100000;
//inst_mem[5]=32'b00000000001000100011000000100010;
//inst_mem[6]=32'b00000000011001000011000000100100;
//inst_mem[7]=32'b00000000001000100011100000100101;
//inst_mem[8]=32'b00000000001000110010100000100110;
//inst_mem[9]=32'b00000000001000100011000000100111;
//inst_mem[10]=32'b00000000100000100011100000000000;
//inst_mem[11]=32'b00000000001000100010100000000010;
//inst_mem[12]=32'b00000000001000010010100000100000;
//inst_mem[13]=32'b00000000101001000011000000100010;
//inst_mem[14]=32'b00000000101001100011100000100100;
//inst_mem[15]=32'b00110100101001010000000000001111;
//inst_mem[16]=32'b10101100000000010000000000000000;
//inst_mem[17]=32'b10101100000001000000000000000100;
//inst_mem[18]=32'b10001100000001010000000000000000;
//inst_mem[19]=32'b10001100000001100000000000000100;
//inst_mem[20]=32'b00110000110001110000000000001011;
//inst_mem[21]=32'b10101100000001110000000000001000;
//inst_mem[22]=32'b10001100000001010000000000000000;
//inst_mem[23]=32'b10101100000001010000000000001100;
//inst_mem[24]=32'b00010000001000010000000000000001;
//inst_mem[25]=32'b00000000010000100010100000100000;
//inst_mem[26]=32'b00010100000000010000000000000010;
//inst_mem[27]=32'b00000000010000100011000000100000;
//inst_mem[28]=32'b00000000100001000011100000100000;
//inst_mem[29]=32'b00001000000000000000000000100000;
//inst_mem[30]=32'b00000000010000100010100000100000;
//inst_mem[31]=32'b00000000100001000011000000100000;
//inst_mem[32]=32'b00000000000000000000000000100000;

	
	
	
	//-------------------------------------------------------------

/* LAST ADDRESS */ inst_mem[2600] = 32'b10110100001000100001100000100000; //Halt 
// every program should end with halt signal 

	

	 
                
            end
            1'b1: begin

          inst_out <= inst_mem[address >> 2];
             
            end
            
        endcase
   
end

endmodule