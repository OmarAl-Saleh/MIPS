module INST_MEM #(
  parameter size = 64,          
  parameter data_width = 32    
)(
 // input clk,
  input reset,                   
  input [31:0] address,
  output reg [31:0] inst_out

);
   reg [31:0] inst_mem [0:size - 1];

  


reg state = 1'b0;
  
  
//  
  always @(*) begin

        case (state)
            1'b0: begin
                state <= 1'b1;
//*******************************************************************************************************


    $readmemh("inst_mem_input.txt", inst_mem);



//*******************************************************************************************************					 
/*
		0- JAL SORT															00001100000000000000000000000010
		1- J   END															00001000000000000000000000011001
SORT	2- LW R16,0(R0)													10001100000100000000000000000000
		3- ADDI R8,R0,R0    //R8=0										00100000000010000000000000000000
		4- ADDI R17,R0,19   //R17=19									00100000000100010000000000010011
SL1	5- BGT  R8,R17,SEL1 //WILL LOOP 19 TIMES					00011001000100010000000000010010 ********************
		6- ADDI R9,R0,0	  //R9=0										00100000000010010000000000000000
		7- SUB  R10,R17,R9   //R10=R17-R9							00000010001010010101000000100010
SL2   8- BGT  R9,R10,SEL2												00011001001010100000000000001101
		9- SLL  R11,R9,2													00000001001000000101100010000000
		10-ADD  R12,R16,R11												00000010000010110110000000100000
		11-LW   R13,0(R12)												10001101100011010000000000000000
		12-LW   R14,4(R12)												10001101100011100000000000000100
		13-BGT  R13,R14,SWAP												00011001101011100000000000000001
		14-J	  ES															00001000000000000000000000010100
SWAP	15-ADD  R15,R13,R0												00000001101000000111100000100000
		16-ADD  R13,R14,R0												00000001110000000110100000100000
		17-ADD  R14,R15,R0												00000001111000000111000000100000
		18-SW   R13,0(R12)												10101101100011010000000000000000
		19-SW   R14,4(R12)												10101101100011100000000000000100
ES		20-ADDI R9,R9,1													00100001001010010000000000000001
		21-J	  SL2															00001000000000000000000000001000
SEL2	22-ADDI R8,R8,1													00100001000010000000000000000001
		23-J	  SL1															00001000000000000000000000000101
SEL1  24-JR	  R31															00000011111001010010000000001000
END	25-ADD R0,R0,R0													00000000000000000000000000100000

LW R1,0(R0)    															10001100000000010000000000000000
LW R2,4(R0)																	10001100000000100000000000000100
LW R3,8(R0)																	10001100000000110000000000001000
LW R4,12(R0)																10001100000001000000000000001100
LW R5,16(R0)																10001100000001010000000000010000
LW R6,20(R0)																10001100000001100000000000010100
LW R7,24(R0)																10001100000001110000000000011000
LW R8,28(R0)																10001100000010000000000000011100
LW R9,32(R0)																10001100000010010000000000100000
LW R10,36(R0)																10001100000010100000000000100100
LW R11,40(R0)																10001100000010110000000000101000
LW R12,44(R0)																10001100000011000000000000101100
LW R13,48(R0)																10001100000011010000000000110000
LW R14,52(R0)																10001100000011100000000000110100
LW R15,56(R0)																10001100000011110000000000111000
LW R16,60(R0)																10001100000100000000000000111100
LW R17,64(R0)																10001100000100010000000001000000
LW R18,68(R0)																10001100000100100000000001000100
LW R19,72(R0)																10001100000100110000000001001000
LW R20,76(R0)																10001100000101000000000001001100
*/

//**********************
/*
10001100000000010000000000000000
00100000000000010000000000000010
10101100000000010000000000000000
10001100000000100000000000000000
*/
//*******************************************************************************************************					 

					 
//		Lw r1,0(R0)		10001100000000010000000000000000				0
//		ori r2 ,r0,4	00110100000000100000000000000100				1
//		addi r3,r0,-2	00100000000000111111111111111110				2
//		Lw r4,4(R0)		10001100000001000000000000000100				3

//		ADD R5,R1,R1	00000000001000010010100000100000				4
//		SUB R6,R1,R2	00000000001000100011000000100010				5
//		AND R6,R3,R4	00000000011001000011000000100100				6
//		OR  R7,R1,R2	00000000001000100011100000100101				7
//		XOR R5,R1,R3	00000000001000110010100000100110				8
//		NOR R6,R1,R2	00000000001000100011000000100111				9
//		SLL R7,R4,R2	00000000100000100011100000000000				10
//		SRL R5,R1,R2	00000000001000100010100000000010				11

//		add r5,r1,r1	00000000001000010010100000100000				12
//		sub r6,r5,r4	00000000101001000011000000100010				13
//		and r7,r5,r6	00000000101001100011100000100100				14
//		ori r5,r5,0xf	00110100101001010000000000001111				15
				
//		sw r1, 0(r0)	10101100000000010000000000000000				16
//		sw r4, 1(r0)	10101100000001000000000000000100				17
//		lw r5, 0(r0)	10001100000001010000000000000000				18
						
//		lw r6,1(r0)		10001100000001100000000000000100				19
//		andi r7,r6,0xb	00110000110001110000000000001011				20
//		sw r7,2(r0)		10101100000001110000000000001000				21
//		lw r5,0(r0)		10001100000001010000000000000000				22
//		sw r5,3(r0)		10101100000001010000000000001100				23


//24           beq r1, r1, P1			00010000001000010000000000000001// 1*4 + 26*4 = 27*4
//             add r5, r2, r2			00000000010000100010100000100000
//P1: 26       bne r0, r1, P2			00010100000000010000000000000010// 2*4 + 28*4 = 30*4
//    27       add r6, r2, r2			00000000010000100011000000100000
//      28     add r7, r4, r4			00000000100001000011100000100000
//P2: 29       j P3						00001000000000000000000000100000
//             add r5, r2, r2			00000000010000100010100000100000
//             add r6, r4, r4			00000000100001000011000000100000
//P3: 32       add r0, r0, r0 		00000000000000000000000000100000



//R1 = F1E0











		
					 // Enter here the Instructions of the program 
					 
					 //*****test for reset *************
		/*			 inst_mem[0] = 32'b10001100000000010000000000000100; //LW R1, 4(R0)
					 inst_mem[1] = 32'b00100000001000010000000000000010; //ADDI R1, R1, 2
					 inst_mem[2] = 32'b10101100000000010000000000000100; //SW R1, 4(R0)
			*/	 
			
			
			
			
	
 /*	inst_mem[0] = 32'b10001100000010000000000000000000; //LW R8, 0(R0)
	inst_mem[1] = 32'b10001100000010010000000000100000; //LW R9, 0x20(R0)
	inst_mem[2] = 32'b10001100000010100000000001010000; //LW R10, 0x50(R0)
	inst_mem[3] = 32'b10001100000010110000000000001000; //LW R11, 0x8(R0)*/
	
	
	/*inst_mem[0] = 32'b10001100000000010000000000000100; //LW R1, 4(R0)      lw r2,56(r0)10001100000000100000000000000000
	inst_mem[1] = 32'b00000000001000100000100010000000; //SLL R1, R1, 2 
	inst_mem[2] = 32'b10101100000000010000000000000100; //SW R1, 4(R0) 
	inst_mem[3] = 32'b10001100000000100000000000010000; //LW R2, 16(R0)
	inst_mem[4] = 32'b10001100000000110000000000010000; //LW R3, 16(R0)
	inst_mem[5] = 32'b00000000010000000001100001000000; //SLL R3, R2, 1 (There is a problem wee need Forwarding to solve it and hazard detection )
	inst_mem[6] = 32'b10101100000000110000000000001100; //SW R3, 12(R0)
	inst_mem[7] = 32'b10001100000001000000000000001100; //LW R4, 12(R0)
*/
	
/*	inst_mem[0] = 32'b00000000000000001110000000000000; //ADD R28,R0,R0 (R28=0)
	inst_mem[1] = 32'b10001111100010000000000000000000; //LW R8, 0(R28)
	inst_mem[2] = 32'b10001111100010010000000000000100; //LW R9, 4(R28)
	inst_mem[3] = 32'b00000001000010010100000000100000; //ADD R8, R8, R9
	inst_mem[4] = 32'b10001111100010100000000000001000; //LW R10, 8(R28)
	inst_mem[5] = 32'b00000001010010100101000000100000; //ADD R10, R10, R10
	inst_mem[6] = 32'b00000001000010100100000000100010; //SUB R8, R8, R10
	inst_mem[7] = 32'b00100001000010000000000000000001; //ADDI R8, R8, 1
	inst_mem[8] = 32'b00000000000010000100000000100010; //SUB R8, R0, R8*/
	
	/*inst_mem[0] = 32'b00000000000000000100000000100000; //ADD R8, R8, R0
	inst_mem[1] = 32'b00100000000010010000000000001010; //ADDI R9, R9, 10
	inst_mem[2] = 32'b00000001000010010101000000100010; //SUB R10, R8, R9 //Loop
	inst_mem[3] = 32'b00100000000011000000000000000001; //ADDI R12, R0, 1
	inst_mem[4] = 32'b00011001000010010000000000000010; //BGT R8, R9, DONE
	inst_mem[5] = 32'b00100001000010000000000000000001; //ADDI R8, R8, 1
	inst_mem[6] = 32'b00001000000000000000000000000010; //JUMP LOOP
	inst_mem[7] = 32'b00000001001000000110100010100000; //ADD R13, R9, R0 //DONE
	inst_mem[8] = 32'b00100000000011100000000000011011; //ADDI R14, R0, 1B(27)
	inst_mem[9] = 32'b00110001110011100000000000010111; //ANDI R14, R14, 17(23)
	*/
	
	/*inst_mem[0] = 32'b00100000000000010000000000000010; //ADDI R1, R0, 2 (a)
	inst_mem[1] = 32'b00100000000000100000000000000010; //ADDI R2, R0, 2 (b)
	inst_mem[2] = 32'b00100000010000110000000000000011; //ADDI R3, R2, 3 (b+3)
	inst_mem[3] = 32'b00100100001000110000000000000010; //BGE  R1, R3, THEN
	inst_mem[4] = 32'b00100000001000010000000000000001; //ADDI R1, R1, 1
	inst_mem[5] = 32'b00001000000000000000000000000111; //JUMP END
	inst_mem[6] = 32'b00100000001000010000000000000010; //ADDI R1, R1, 2 //THEN 
	inst_mem[7] = 32'b00000000010000010001000000100000; //ADD R2, R2, R1 //END*/
	
	/*inst_mem[0] = 32'b00100000000000010000000000000110; //ADDI R1, R0, 6 (a)
	inst_mem[1] = 32'b00100000000000100000000000000010; //ADDI R2, R0, 2 (b)
	inst_mem[2] = 32'b00100000010000110000000000000011; //ADDI R3, R2, 3 (b+3)
	inst_mem[3] = 32'b00100100001000110000000000000010; //BGE  R1, R3, THEN
	inst_mem[4] = 32'b00100000001000010000000000000001; //ADDI R1, R1, 1
	inst_mem[5] = 32'b00001000000000000000000000000111; //JUMP END
	inst_mem[6] = 32'b00100000001000010000000000000010; //ADDI R1, R1, 2 //THEN 
	inst_mem[7] = 32'b00000000010000010001000000100000; //ADD R2, R2, R1 //END*/
	
	/*inst_mem[0] = 32'b00000000000000000000100000100000; //ADD R1, R0, R0 
	inst_mem[1] = 32'b00000000000000000001000000100000; //ADD R2, R0, R0
	inst_mem[2] = 32'b00100000000010010000000001100100; //ADDI R9, R0, 100
	inst_mem[3] = 32'b00010000001010010000000000000010; //BEQ R1, R9, EXIT //START
	inst_mem[4] = 32'b00100000001000010000000000000001; //ADDI R1, R1, 1
	inst_mem[5] = 32'b00001000000000000000000000000011; //JUMP START
	inst_mem[6] = 32'b00000000001000100001100000100000; //ADD R3, R0, R0 //EXIT*/
	
	
//-------------------------------------------------------------

//

/* LAST ADDRESS */ //inst_mem[3] = 32'b10110100001000100001100000100000; //Halt B4221820
// every program should end with halt signal 

	/*
	BENCHMARK1
	
8C010000
34020004
2003FFFE
8C040004
00212820
00223022
00643024
00223825
00232826
00223027
00823800
00222802
00212820
00A43022
00A63824
34A5000F
AC010000
AC040004
8C050000
8C060004
30C7000B
AC070008
8C0A0000
AC05000C
10210001
00422820
14010002
00423020
00843820
08000020
00422820
00843020
00000020
B4221820
	
	
	*/
	
	/*
	
	BM2
	0C000002
08000019
8C100000
20080000
20110013
19110012
20090000
02295022
192A000D
01205880
020B6020
8D8D0000
8D8E0004
19AE0001
08000014
01A07820
01C06820
01E07020
AD8D0000
AD8E0004
21290001
08000008
21080001
08000005
03E00008
00000020
B4221820
	*/

	 
                
            end
            1'b1: begin
	
          inst_out <= inst_mem[address >> 2];
            end

        endcase
    end
//end

endmodule